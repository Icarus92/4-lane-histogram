library verilog;
use verilog.vl_types.all;
entity histogram_lane_tb is
end histogram_lane_tb;
